module fulladder(input logic a, b, cin,
                   output logic s, cout);

  logic p, g;
  always_comb
  begin
    p = a ^ b; // blocking
    g = a & b; // blocking
    s = p ^ cin; // blocking
    cout = g | (p & cin); // blocking
  end
  
endmodule
